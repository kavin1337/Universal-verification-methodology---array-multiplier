interface mul_interface();
  
  logic [3:0] a,b;
  logic [7:0] p;
  
  
endinterface: mul_interface
